module or_gate(
				input wire d,e,
				output wire f
				);
				
				
				assign f = d | e;
				
				
endmodule
